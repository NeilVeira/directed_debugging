../../sva/wb_dma_inc30r.sv