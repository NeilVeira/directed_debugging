../../sva/wb_dma_ch_rf.sv