../../sva/wb_dma_wb_if.sv