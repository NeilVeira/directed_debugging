../../../tb/include/sel_test.vh