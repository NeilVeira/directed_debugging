../../sva/wb_dma_de.sv