../../sva/wb_dma_top.sv