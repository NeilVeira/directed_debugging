../../sva/except.sv