../../sva/wb_dma_ch_arb.sv