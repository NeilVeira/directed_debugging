../../sva/wb_dma_ch_pri_enc.sv