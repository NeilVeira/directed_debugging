../../../sva/include/func.sv