../../sva/fpu.sv