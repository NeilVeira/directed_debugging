../../sva/pre_norm.sv