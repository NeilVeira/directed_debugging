../../sva/wb_dma_ch_sel.sv