../../sva/post_norm.sv