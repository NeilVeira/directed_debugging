../../sva/wb_dma_rf.sv