../../sva/assumption.sv